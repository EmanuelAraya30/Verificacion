module compuerta (E1,E2,S1);

	input E1, E2;
	output S1;

	assign S1 = E1 & E2;

endmodule
